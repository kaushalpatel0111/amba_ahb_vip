// AHB Package
`ifndef AHB_PKG
`define AHB_PKG

`include "ahb_top_define.svh"
`include "ahb_topvar_define.sv"
`include "ahb_mas_intf.sv"
`include "ahb_slv_intf.sv"
//`include "ahb_common_intf.sv"
`include "ahb_checker.sv"

package ahb_pkg;
    // uvm
     import uvm_pkg::*;
    `include "uvm_macros.svh"

    // define
    `include "ahb_top_define.svh"
    `include "ahb_topvar_define.sv"
    `include "ahb_enum_pkg.sv"

    // config
    `include "ahb_cfg.sv"
    `include "ahb_mas_cfg.sv"
    `include "ahb_slv_cfg.sv"
    `include "ahb_sys_cfg.sv"
    `include "ahb_cust_cfg.sv"

    // ahb base transaction
    `include "ahb_transaction.sv"	

    // ahb memory
    `include "ahb_slv_mem.sv"

    // sequence
    `include "ahb_base_seq.sv"
    
    // ahb master
    `include "ahb_mas_seq_item.sv"
    `include "ahb_mas_base_seq.sv"
    `include "ahb_mas_single_burst_trans_seq.sv"
    `include "ahb_mas_incr4_burst_trans_seq.sv"
    `include "ahb_mas_incr_undefined_len_burst_trans_seq.sv"
    `include "ahb_mas_incr8_burst_trans_seq.sv"
    `include "ahb_mas_incr16_burst_trans_seq.sv"
    `include "ahb_mas_wrap4_burst_trans_seq.sv"
    `include "ahb_mas_wrap8_burst_trans_seq.sv"
    `include "ahb_mas_wrap16_burst_trans_seq.sv"
    `include "ahb_mas_busy_during_fixed_burst_trans_seq.sv"
    `include "ahb_mas_narrow_trans_seq.sv"
    `include "ahb_mas_error_seq.sv"
    `include "ahb_mas_random_burst_seq.sv"
    `include "ahb_mas_seqr.sv"
    `include "ahb_mas_drv.sv"
    `include "ahb_mas_mon.sv"
    `include "ahb_mas_agnt.sv"

    // ahb slave
    `include "ahb_slv_seq_item.sv"
    `include "ahb_slv_seqr.sv"
    `include "ahb_slv_base_seq.sv"
    `include "ahb_slv_drv.sv"
    `include "ahb_slv_mon.sv"
    `include "ahb_slv_agnt.sv"

    // reset sequence
    `include "ahb_rst_seq.sv"

    // env
    `include "ahb_mas_fc.sv"
    `include "ahb_slv_fc.sv"
    `include "ahb_scb.sv"
    `include "ahb_env.sv" 

    // base test
    `include "ahb_base_test.sv"

    // testcases
    `include "ahb_sanity_test.sv"
    `include "ahb_in_bw_rst_test.sv"
    `include "ahb_single_burst_trans_test.sv"
    `include "ahb_incr_undefined_len_burst_trans_test.sv"
    `include "ahb_incr4_burst_trans_test.sv"
    `include "ahb_incr8_burst_trans_test.sv"
    `include "ahb_incr16_burst_trans_test.sv"    
    `include "ahb_wrap4_burst_trans_test.sv"    
    `include "ahb_wrap8_burst_trans_test.sv"    
    `include "ahb_wrap16_burst_trans_test.sv"    
    `include "ahb_busy_during_fixed_burst_trans_test.sv"    
    `include "ahb_busy_during_undefined_len_burst_trans_test.sv"    
    `include "ahb_narrow_trans_test.sv"    
    `include "ahb_error_injection_test.sv"    
    `include "ahb_random_burst_trans_test.sv"    
    
endpackage

`endif
