// AHB TOP Define
`ifndef AHB5
	`define AHB5
`endif
