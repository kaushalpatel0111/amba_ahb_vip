// AHB Base Test 
`ifndef AHB_BASE_TEST
`define AHB_BASE_TEST

class ahb_base_test extends uvm_test;
    
    `uvm_component_utils(ahb_base_test)

    ahb_cust_cfg cust_cfg_h;
    ahb_env env_h;
    
    function new(string name = "ahb_base_test", uvm_component parent = null);
        super.new(name, parent);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
      
      	cust_cfg_h = ahb_cust_cfg::type_id::create("cust_cfg_h", this);
      	
      	if (!uvm_config_db #(virtual ahb_mas_intf)::get(this,"env_h.magnt_h", "ahb_mas_intf", cust_cfg_h.mcfg_h.mvif))
          `uvm_fatal("MINTF_FATAL", "Configuration object of Master vif is not set properly");
      
        if (!uvm_config_db #(virtual ahb_slv_intf)::get(this,"env_h.sagnt_h", "ahb_slv_intf", cust_cfg_h.scfg_h.svif))
          `uvm_fatal("SINTF_FATAL", "Configuration object of Slave vif is not set properly");
      
      	env_h = ahb_env::type_id::create("env_h", this);
        
	//set cust configure
        uvm_config_db #(ahb_cust_cfg)::set(this,"*", "ahb_cust_cfg", cust_cfg_h);
    endfunction

    function void end_of_elaboration_phase(uvm_phase phase);
      	//cust_cfg_h.print();
    endfunction

    function void report_phase(uvm_phase phase);
        uvm_report_server svr_h;

        //is a global server that processes all of the reports generated by a uvm_report_handler.
        //get server method of uvm report server return get_report_server  

        svr_h = uvm_report_server::get_server();

        if((svr_h.get_severity_count(UVM_WARNING) + svr_h.get_severity_count(UVM_FATAL) + svr_h.get_severity_count(UVM_ERROR)) == 0)begin
            `uvm_info("REPORT PHASE","TEST PASS !!",UVM_NONE)
            // method are get_severity return number of counts of uvm_fatal,warning,error
            $display("");
            $display("  ######  ######  ######  ###### ");
            $display("  #    #  #    #  #       #     ");
            $display("  #    #  #    #  #       #     ");
            $display("  #    #  #    #  #       #     ");
            $display("  ######  ######  ######  ###### ");
            $display("  #       #    #       #       # ");
            $display("  #       #    #       #       # ");
            $display("  #       #    #       #       # ");
            $display("  #       #    #  ######  ###### ");
            $display("");

        end
        else begin
            `uvm_info("REPORT PHASE","TEST FAIL !!",UVM_NONE)
            
            $display("");
            $display("  ######  ######  #######  #      ");
            $display("  #       #    #     #     #      ");
            $display("  #       #    #     #     #      ");
            $display("  #       #    #     #     #      ");
            $display("  ######  ######     #     #      ");
            $display("  #       #    #     #     #      ");
            $display("  #       #    #     #     #      ");
            $display("  #       #    #     #     #      ");
            $display("  #       #    #  #######  ####### ");
            $display("");
            
            //$finish;

        end
    endfunction

endclass

`endif
